--
-- Copyright (c) 2023 Charlie Amtorp
--
-- Permission is hereby granted, free of charge, to any person
-- obtaining a copy of this software and associated documentation
-- files (the "Software"), to deal in the Software without
-- restriction, including without limitation the rights to use,
-- copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the
-- Software is furnished to do so, subject to the following
-- conditions:
--
-- The above copyright notice and this permission notice shall be
-- included in all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
-- EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
-- OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
-- NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
-- HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
-- WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
-- OTHER DEALINGS IN THE SOFTWARE.
--

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
	use ieee.std_logic_unsigned.all;

use work.CoreTypes.all;

entity AluShiftBlock is

	port
	(
		InstSWAP	: in  std_logic;
		InstLSR		: in  std_logic;
		InstASR		: in  std_logic;
		InstROR		: in  std_logic;
		
        A			: in  DataWord;
        iC			: in  std_logic;                   
		
		oV			: out std_logic;
		oC			: out std_logic;
		result		: out DataWord
	);
	
end entity;
	
architecture RTL of AluShiftBlock is

	signal tmp : DataWord;

begin
	result <= tmp;

	SFT : process(InstSWAP, InstLSR, InstASR, InstROR, A, iC) begin
	
		tmp(3 downto 0) <= A(7 downto 4);
		tmp(7 downto 4) <= A(3 downto 0);
		oV <= '0';
		oC <= '0';

		if InstLSR then
	
			tmp(7) <= '0';
			tmp(6 downto 0) <= A(7 downto 1);
			oC <= A(0);
			oV <= A(0) xor '0';
			
		elsif InstASR then
	
			tmp(7) <= A(7);
			tmp(6 downto 0) <= A(7 downto 1);
			oC <= A(0);
			oV <= A(0) xor A(7);
			
		elsif InstROR then
			
			tmp(7) <= iC;
			tmp(6 downto 0) <= A(7 downto 1);
			oC <= A(0);
			oV <= A(0) xor iC;
			
		end if;
	
	end process;
	
end architecture;