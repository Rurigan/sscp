--
-- Copyright (c) 2023 Charlie Amtorp
--
-- Permission is hereby granted, free of charge, to any person
-- obtaining a copy of this software and associated documentation
-- files (the "Software"), to deal in the Software without
-- restriction, including without limitation the rights to use,
-- copy, modify, merge, publish, distribute, sublicense, and/or sell
-- copies of the Software, and to permit persons to whom the
-- Software is furnished to do so, subject to the following
-- conditions:
--
-- The above copyright notice and this permission notice shall be
-- included in all copies or substantial portions of the Software.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
-- EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES
-- OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
-- NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT
-- HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY,
-- WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
-- OTHER DEALINGS IN THE SOFTWARE.
--

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;
	use ieee.std_logic_unsigned.all;

use work.CoreTypes.all;

entity ProcessorMemory is

	generic 
	(
		ProgramFile : string := "(none)"
	);

	port
	(
		SysCtrl			: in	SystemCtrlRec;
		ToPrgMem		: in 	PrgMemoryCtrlRec;
		ToDataMem		: in 	DataMemoryCtrlRec;
		FromPrgMem		: out	PrgMemoryOutRec;
		FromDataMem		: out 	DataMemoryOutRec
	);

end entity;

architecture RTL of ProcessorMemory is

begin

	PRG : component ProgramMemory 

		generic map
		(
			InitFile 	=>	ProgramFile
		)

		port map 
		(
			SysCtrl		=>	SysCtrl,
			FromCpu		=>	ToPrgMem,
			ToCpu		=>	FromPrgMem
		);
		
		
	DATA : component DataMemory

		port map
		(
			SysCtrl		=>	SysCtrl,
			FromCpu		=>	ToDataMem,
			ToCpu		=>	FromDataMem
		);

end architecture;